module mult4_4
(
input [3:0]data_a,
input [3:0]data_b,
output[7:0]product_
);
assign product_ = data_a * data_b;
endmodule
